module fpga_top;
    // Temporary stub top module
endmodule
